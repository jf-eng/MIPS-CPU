module regfile (
	
);
	

	
endmodule