module ram (
	ports
);
	
endmodule