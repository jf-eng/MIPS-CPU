module rom (
	ports
);
	
endmodule