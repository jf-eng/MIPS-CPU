module datapath (
	ports
);
	
endmodule