module regfile_tb ();
	
	regfile dut();


endmodule