module alu(
	input logic[31:0] op1, op2,
	input logic Add, Sub, Mul, Div, Unsigned, 
	input Or, And, Xor, SL, SR, Arithmetic,
	output logic[31:0] alu_out
);


endmodule