module controlpath (
	ports
);
	
endmodule